parameter DIN_WIDTH=16;
parameter M=2;
parameter N=4;
parameter R=500;
parameter DOUT_WIDTH=56;
parameter MODE=0;
