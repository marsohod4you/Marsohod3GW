parameter DIN_WIDTH = 16;
parameter COEFF_WIDTH = 16;
parameter DOUT_WIDTH = 31;
parameter NUM_CHN = 2;
parameter NUM_FACTOR = 2;
parameter TAPS_SIZE = 23;
parameter NUM_TDM = 1;
parameter COEFF_PATH = "./coeff.dat";
