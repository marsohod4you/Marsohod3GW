`define MODULE_NAME CIC_Fliter_Top
`define DECIMATOR
